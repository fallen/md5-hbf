module top(input clock, input reset, output led, output led2, output led3);

generator g1 (clock, reset, led);

endmodule
